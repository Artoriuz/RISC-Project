library verilog;
use verilog.vl_types.all;
entity memtest_vlg_vec_tst is
end memtest_vlg_vec_tst;
