library verilog;
use verilog.vl_types.all;
entity microprocessador_vlg_vec_tst is
end microprocessador_vlg_vec_tst;
